module main

import graphics

fn main() {
	mut app := graphics.create_app()
	graphics.run(mut app)
}
