module egg

import ecs

pub struct IsEggTag {
	ecs.ComponentBase
}
