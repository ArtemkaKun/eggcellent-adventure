module common

import transform

pub struct Entity {
pub:
	position transform.Position
	image_id int
}
