module common

// Orientation represents the direction an object is facing or moving in the game world.
// used for rendering and calculations.
pub enum Orientation {
	left
	right
}
