module main

import graphics

fn main() {
	mut app := graphics.create_app()
	graphics.start_app(mut app)
}
