module world

import obstacle

pub struct Model {
pub:
	obstacle_positions []obstacle.Position
}
